package timing_constants_tb;

  // Timing constants in nanoseconds for simulation
  localparam time T1H_NS = 700;  // 700 ns
  localparam time T1L_NS = 600;  // 600 ns
  localparam time T0H_NS = 350;  // 350 ns
  localparam time T0L_NS = 800;  // 800 ns
  localparam time TRESET_NS = 50000;  // Reset duration (50 µs)

endpackage
