/*
-----------------------------------------------------------------------------
Module Name: timer
Description: Encapsulates the count_enable and counter modules.

Author: Curtis Button
Date: March 19, 2025
-----------------------------------------------------------------------------
*/

`include "count_enable.sv"
`include "counter.sv"

module timer (
    input logic i_clk,          // Clock input
    input logic i_reset_n,      // Active low reset
    input logic i_rising,       // Synchronized rising edge for LED control
    input logic i_falling,      // Synchronized falling edge for LED control
    output pipeline_types::decoder_input_t#(10) o_count // Counter output signal
);

    //////////////////////////////////////////////////////////////////////
    // Internal Signals
    logic w_count_enable;  // Clock enable signal generated by count_enable

    //////////////////////////////////////////////////////////////////////
    // Instance: Count Enable
    // Generates a clock enable signal by dividing the input clock
    count_enable u_count_enable (
        .i_clk(i_clk),
        .i_reset_n(i_reset_n),
        .i_rising(i_rising),
        .o_count_enable(w_count_enable)
    );

    //////////////////////////////////////////////////////////////////////
    // Instance: Counter
    // Increments the counter based on the clock enable signal
    counter u_counter (
        .i_clk(i_clk),
        .i_reset_n(i_reset_n),
        .i_count_enable(w_count_enable),
        .i_rising(i_rising),
        .i_falling(i_falling),
        .o_count(o_count)
    );

endmodule