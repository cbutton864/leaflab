interface led_if;
  logic serial_in;
  logic [23:0] o_led_data;
  logic rst_n;
endinterface
